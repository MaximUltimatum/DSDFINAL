`timescale 1ns / 1ps

module toggle_motor(
    input  rf_in,
    input  sw_in,
    output out
    );
    
    wire rf_db_in;
    wire sw_in;

endmodule
