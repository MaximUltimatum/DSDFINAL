`timescale 1ns / 1ps

module toggle_lock(
    input in,
    output out
    );

endmodule
