`timescale 1ns / 1ps

module rf_controller(

    );



endmodule
