`timescale 1ns / 1ps

module debouce(

    );


endmodule
