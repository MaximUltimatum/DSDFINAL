`timescale 1ns / 1ps

module toggle_motor(
    input  rf_in,
    input  sw_in,
    output out
    );

endmodule
